`default_nettype none
module quick_uart_rx #(
    parameter BAUD = 115200,
    parameter DATA_BITS = 8,
    parameter STOP_BITS = 1,
) (
);
endmodule
`default_nettype wire

